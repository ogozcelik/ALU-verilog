//TESTBENCH

`timescale 1ns/1ps
module ALU_design_tb();

reg clk;
reg [31:0] A,B;
reg [4:0] ALU_CONTROL;
wire [31:0] Y;
wire Z, V, N, C;

// instantiate device under test
ALU_design dut(A,B,ALU_CONTROL,clk,Y,Z, V, N, C);

always begin
	clk = 0; #5; clk = 1; #5;
end

initial begin
//addition check
A = 32'b10000000000000000000000000010000; B=32'b00000000000000000000000000000100; ALU_CONTROL=5'b00000; #20; // -16 + 4 = -12
if (Y !== 32'b10000000000000000000000000001100) $display ("addition failed.");
if (Z !== 0 && V !== 0 && N !== 1 && C !== 0) $display ("flags failed.");

//subtraction check
A = 32'b00000000000000000000000001010010; B=32'b00000000000000000000000000100000; ALU_CONTROL=5'b00001; #20; // 82 - 32 = 50
if (Y !== 32'b00000000000000000000000000110010) $display ("subtraction failed.");
if (Z !== 0 && V !== 0 && N !== 0 && C !== 0) $display ("flags failed.");

//multiplication check
A = 32'b00000000000000001000000000000010; B=32'b00000000000000000000000000000111; ALU_CONTROL=5'b00010; #20; // -2 * 7 = -14
if (Y !== 32'b10000000000000000000000000001110) $display ("multiplication failed.");
if (Z !== 0 && V !== 0 && N !== 1 && C !== 0) $display ("flags failed.");

//divison check
A = 32'b00000000000000000000000000010111; B=32'b00000000000000000000000000000110; ALU_CONTROL=5'b00011; #20; // 23 / 6 = quot 3, remainder 5
if (Y !== 32'b00000000000000101000000000000011) $display ("division failed.");
if (Z !== 0 && V !== 0 && N !== 0 && C !== 0) $display ("flags failed.");

//bit-wise and
A = 32'b01000010000110000000001100000010; B=32'b10111101111001111111110011111101; ALU_CONTROL=5'b01000; #20;
if (Y !== 32'b00000000000000000000000000000000) $display ("bw and failed.");

//bit-wise or
A = 32'b01000010000110000000001100000010; B=32'b00000000000000000000000000000000; ALU_CONTROL=5'b01001; #20;
if (Y !== 32'b01000010000110000000001100000010) $display ("bw or failed.");

//bit-wise xor
A = 32'b00000010010100000001100000000010; B=32'b00000010000100000001100000000000; ALU_CONTROL=5'b01010; #20;
if (Y !== 32'b00000000010000000000000000000010) $display ("bw xor failed.");

//bit-wise nor
A = 32'b11111000000000000000000000000010; B=32'b00000000000000000000000000000000; ALU_CONTROL=5'b01011; #20;
if (Y !== 32'b00000111111111111111111111111101) $display ("bw nor failed.");

//bit-wise nand
A = 32'b10000000000000000000000000111000; B=32'b10000000000000000000000000111000; ALU_CONTROL=5'b01100; #20;
if (Y !== 32'b01111111111111111111111111000111) $display ("bw nand failed.");

//bit-wise xnor
A = 32'b01010100000000000000000000000000; B=32'b01010101111111111111111100000000; ALU_CONTROL=5'b01101; #20;
if (Y !== 32'b11111110000000000000000011111111) $display ("bw xnor failed.");

//compare EQ
A = 32'b10000000000000000000000000000000; B=32'b00000000000000000000000000000000; ALU_CONTROL=5'b10000; #20; // check a special case where -0 ?== +0
if (Y !== 32'b00000000000000000000000000000001) $display ("compare eq 1 failed.");

//compare EQ
A = 32'b10000000000000000000000000011000; B=32'b10000000000000000000000000011000; ALU_CONTROL=5'b10000; #20; // -24 ?== -24 => yes
if (Y !== 32'b00000000000000000000000000000001) $display ("compare eq 2 failed.");

//compare LT
A = 32'b10000000000000000000000000110000; B=32'b00000000000000000000000000000100; ALU_CONTROL=5'b10001; #20; // -48 ?< +4 => yes
if (Y !== 32'b00000000000000000000000000000010) $display ("compare lt failed.");

//COMPARE GT
A = 32'b10000000000000000000000000000010; B=32'b10000000000000000000000000100001; ALU_CONTROL=5'b10010; #20; // -2 ?> -33 => yes
if (Y !== 32'b00000000000000000000000000000100) $display ("compare gt failed.");

//LSL
A = 32'b11000000000000000000000001101110; B=32'b00000000000000000000000000000010; ALU_CONTROL=5'b11000; #20; // 2 bit lsl
if (Y !== 32'b00000000000000000000000110111000) $display ("LSL failed.");

//LSR	
A = 32'b10100000000000000000000001101110; B=32'b00000000000000000000000000000011; ALU_CONTROL=5'b11001; #20; // 3 bit lsr
if (Y !== 32'b00010100000000000000000000001101) $display ("LSR failed.");

//ASR
A = 32'b10000000000000000000010111101010; B=32'b00000000000000000000000000001000; ALU_CONTROL=5'b11010; #20; // 8 bit asr
if (Y !== 32'b11111111100000000000000000000101) $display ("ASR failed.");

//REV
A = 32'b10000000000000000000000011000110; ALU_CONTROL=5'b11011; #50;
if (Y !== 32'b01100011000000000000000000000001) $display ("REV failed.");

$display ("END OF TESTBENCH / OGUZHAN OZCELIK 2232544");
$display ("There might be red lines for the outputs for a 15ns since I did not give any initial value to them!");
end


endmodule
